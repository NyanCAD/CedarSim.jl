// Simplified SkyWater nfet_01v8 model (single bin from w=1e-6, l=0.5e-6)

parameters sky130_fd_pr__nfet_01v8__toxe_slope_spectre=0.0
parameters sky130_fd_pr__nfet_01v8__vth0_slope_spectre=0.0
parameters sky130_fd_pr__nfet_01v8__voff_slope_spectre=0.0

subckt sky130_fd_pr__nfet_01v8 (d g s b)
parameters l=1 w=1 nf=1.0 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1
msky130_fd_pr__nfet_01v8 (d g s b) sky130_fd_pr__nfet_01v8__model l=l w=w nf=nf ad=ad as=as pd=pd ps=ps nrd=nrd nrs=nrs sa=sa sb=sb sd=sd
ends

// Load BS IM4 device model
load "spice/bsim4v8.osdi"

// Model for w=1.0e-6, l=0.5e-6  (falls in bin: 4.2e-7 < w < 5.2e-7, 1.5e-7 < l < 1.8e-7)
model sky130_fd_pr__nfet_01v8__model sp_bsim4v8 ( type=1 lmin=1.5e-07 lmax=1.8e-07 wmin=4.2e-07 wmax=5.2e-7 toxe=4.148e-09 toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0=1.442666050e+00 lvth0=-1.228100366e-07 wvth0=-3.135030950e-07 pvth0=3.652871475e-14 k1=0.90707349 k2=-5.135550875e-03 lk2=-1.458596362e-08 wk2=-6.049227457e-08 pk2=6.808591163e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-7.653070645e-01 ldsub=9.410246186e-08 wdsub=5.226696447e-07 pdsub=-3.540906255e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000005e-03 lcdscd=-6.359062582e-19 wcdscd=-1.896999918e-18 pcdscd=2.392799500e-25 cit=0.0 voff=-2.075300007e-01 lvoff=8.330447443e-17 wvoff=2.485092132e-16 pvoff=-3.134598137e-23 nfactor=2.562288561e+01 lnfactor=-2.784724284e-06 wnfactor=-1.126386412e-05 pnfactor=1.363601460e-12 eta0=-1.136614502e-02 leta0=1.774664763e-09 weta0=4.276876208e-09 peta0=-6.677744065e-16 etab=-0.043998 u0=1.518526513e-01 lu0=-1.640557596e-08 wu0=-5.918769347e-08 pu0=7.923070781e-15 ua=-1.793883530e-09 lua=8.618821411e-17 wua=2.903304318e-16 pua=-4.081658001e-23 ub=8.336513898e-18 lub=-9.440161977e-25 wub=-3.672387679e-24 pub=5.526257949e-31 uc=-4.845095256e-10 luc=7.917999472e-17 wuc=2.534405742e-16 puc=-3.552638160e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.951236289e+05 lvsat=-1.568267986e-02 wvsat=-5.697714417e-02 pvsat=8.256077967e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.261698858e-02 lketa=2.206317671e-08 wketa=1.702702291e-08 pketa=-1.423641446e-14 dwg=0.0 dwb=0.0 pclm=-2.686070209e-02 lpclm=3.115085549e-08 wpclm=1.374092151e-07 ppclm=-2.095516005e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-3.930083952e-07 lalpha0=5.335658687e-14 walpha0=2.014712848e-13 palpha0=-2.541278195e-20 alpha1=0.85 beta0=3.404518278e+00 lbeta0=1.317551282e-06 wbeta0=5.007551470e-06 pbeta0=-6.316325119e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-4.010308949e-01 lkt1=2.019060909e-08 wkt1=9.939896227e-08 pkt1=-1.253778751e-14 kt2=-0.028878939 at=2.495577075e+05 lat=-2.470212364e-02 wat=-9.327374313e-02 pat=1.176517686e-8 ute=-1.851973592e+00 lute=6.215089330e-08 wute=1.206579809e-07 pute=-8.564988193e-15 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0 )
